module bist_controller(
    input wire start,
    input wire rst,
    input wire clk,
    output wire test_mode,
    output wire dut_start,
    output wire crc_start,
    output reg[7:0] a_lfsr,
    output reg[7:0] b_lfsr,
    output reg[7:0] test_mode_ctr
);
    

endmodule
