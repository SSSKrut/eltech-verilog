module bist_controller(
    input wire test,
    output wire bist_test,
    output reg[7:0] a_lfsr,
    output reg[7:0] b_lfsr,
    output reg[7:0] bist_out
);
    

endmodule
