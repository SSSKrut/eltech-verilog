module crc8 (
    input reg[7:0] y_in,
    input wire start,
    input wire rst,
    input wire clk,
    output reg[7:0] crc_result
);

endmodule